library verilog;
use verilog.vl_types.all;
entity tutorial_1_vlg_vec_tst is
end tutorial_1_vlg_vec_tst;
